 * @Author: Donald duck tang5722917@163.com
 * @Date: 2023-06-21 15:31:10
 * @LastEditors: Donald duck tang5722917@163.com
 * @LastEditTime: 2023-06-21 15:32:37
 * @FilePath: \spice_netlist_front_end\test\Base\05_ISource_two_resistor\05_ISource_two_resistor.cir
 * @Description: 1 Current Source and two resistor
 * Copyright (c) 2023 by Donald duck email: tang5722917@163.com, All Rights Reserved.
 */

I1 0 1 DC 1A
R1 1 2 1ohm
R2 2 0 3.3ohm 
.OP

.control
    set filetype = ascii
.endc
.end
